// uvm_classic/sequencers/cpu_instruction_sequencer.sv
//
// Copyright (c) 2025 Igor Bogdanov
// All rights reserved.

typedef uvm_sequencer#(riscv_instruction_transaction) cpu_instruction_sequencer; 